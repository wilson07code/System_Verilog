package my_package;

typedef enum{red,green,blue}colors;

typedef struct{

int field_a;
colors c;
}mystruct;

endpackage